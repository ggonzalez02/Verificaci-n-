module Adder (
    input Signo,
    input [7:0] Exp_comun,
    input [25:0] Resul_Mantissa_A,
    input [25:0] Resul_Mantissa_B,
    output[23:0] Suma_resul
);
    
endmodule