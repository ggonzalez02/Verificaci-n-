//////////////////////////////////////////////////////////////////////////////////
// University:  Instituto Tecnológico de Costa Rica                             
// Engineers:   Anthony Artavia                                                 
//              Maricruz Campos                                                 
//              Gabriel González                                                
//  
// Module Name: queue
// Description: 
//////////////////////////////////////////////////////////////////////////////////
module queue (input EN, input CLK, input RST,);
input  [7:0] DATA ;
output [31:0] Data_Q;
wire a, b , c ;






endmodule 