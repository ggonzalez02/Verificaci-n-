//////////////////////////////////////////////////////////////////////////////////
// University:  Instituto Tecnológico de Costa Rica                             
// Engineers:   Anthony Artavia                                                 
//              Maricruz Campos                                                 
//              Gabriel González                                                
//  
// Module Name: Registros
// Description:
//////////////////////////////////////////////////////////////////////////////////
module registros88 (input clk, input rst, input data, );




endmodule  