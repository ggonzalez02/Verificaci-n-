//////////////////////////////////////////////////////////////////////////////////
// University:  Instituto Tecnológico de Costa Rica                             
// Engineers:   Anthony Artavia                                                 
//              Maricruz Campos                                                 
//              Gabriel González                                                
//  
// Module Name: top
// Description: Módulo top de la interfaz
//////////////////////////////////////////////////////////////////////////////////

module top (
    input clk,
    input reset,
    input [2:0] OP,
    input [2:0] Reg1,
    input [2:0] Reg2,
    inout RD_WR,
    inout [7:0] Data,
    output [19:0] Direction
);
    //Definicion de señales internas

    //Banco de registros

    //Segmentos

    //Queue

    //ALU

    
endmodule