//////////////////////////////////////////////////////////////////////////////////
// University:  Instituto Tecnológico de Costa Rica                             
// Engineers:   Anthony Artavia                                                 
//              Maricruz Campos                                                 
//              Gabriel González                                                
//  
// Module Name: queue
// Description: 
//////////////////////////////////////////////////////////////////////////////////
module queue (
    input EN;
    input clk;
    input rst;
    input  [7:0] data ;
    output [31:0] Data_Q;
);

// Data -> R1 -> R2 -> R3 -> R4
wire [7:0] OUT1,OUT2,OUT3,OUT4 

reg





endmodule 