//////////////////////////////////////////////////////////////////////////////////
// University:  Instituto Tecnológico de Costa Rica                             
// Engineers:   Anthony Artavia                                                 
//              Maricruz Campos                                                 
//              Gabriel González                                                
//  
// Module Name: Regsitros de Segmentos
// Description:
//////////////////////////////////////////////////////////////////////////////////

module segments (
    input wire clk;
    input wire rst; 
    output [15:0] segmento;
);




endmodule
