module Desnormalizador (
    input  [23:0] Mantissa_A,
    input  [7:0]  Exponente_A,
    input  [23:0] Mantissa_B,
    input  [23:0] Exponente_B,
    output [25:0] Resul_Mantissa_A,
    output [7:0]  Exp_comun,
    output [23:0] Resul_Mantissa_B
);
// Alinear Mantissa 

// Sacar resultado de exponente comun si ambos exponentes son diferentes 


endmodule