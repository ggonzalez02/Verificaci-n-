module Normalizador (
    input OP_input,
    input Signo,
    input [7:0]  Exp_resul,
    input [47:0] Producto,
    input [25:0] Suma_resul, 
    output[31:0] Resultado
);
    
endmodule